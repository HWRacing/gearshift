// ADCTestADC.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module ADCTestADC (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         altpll_0_c0_clk;                                            // altpll_0:c0 -> modular_adc_0:adc_pll_clock_clk
	wire         altpll_0_locked_conduit_export;                             // altpll_0:locked -> modular_adc_0:adc_pll_locked_export
	wire  [31:0] master_0_master_readdata;                                   // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                                // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                    // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                       // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                 // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                              // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                      // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                  // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire  [31:0] mm_interconnect_0_modular_adc_0_sample_store_csr_readdata;  // modular_adc_0:sample_store_csr_readdata -> mm_interconnect_0:modular_adc_0_sample_store_csr_readdata
	wire   [6:0] mm_interconnect_0_modular_adc_0_sample_store_csr_address;   // mm_interconnect_0:modular_adc_0_sample_store_csr_address -> modular_adc_0:sample_store_csr_address
	wire         mm_interconnect_0_modular_adc_0_sample_store_csr_read;      // mm_interconnect_0:modular_adc_0_sample_store_csr_read -> modular_adc_0:sample_store_csr_read
	wire         mm_interconnect_0_modular_adc_0_sample_store_csr_write;     // mm_interconnect_0:modular_adc_0_sample_store_csr_write -> modular_adc_0:sample_store_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_0_sample_store_csr_writedata; // mm_interconnect_0:modular_adc_0_sample_store_csr_writedata -> modular_adc_0:sample_store_csr_writedata
	wire  [31:0] mm_interconnect_0_modular_adc_0_sequencer_csr_readdata;     // modular_adc_0:sequencer_csr_readdata -> mm_interconnect_0:modular_adc_0_sequencer_csr_readdata
	wire   [0:0] mm_interconnect_0_modular_adc_0_sequencer_csr_address;      // mm_interconnect_0:modular_adc_0_sequencer_csr_address -> modular_adc_0:sequencer_csr_address
	wire         mm_interconnect_0_modular_adc_0_sequencer_csr_read;         // mm_interconnect_0:modular_adc_0_sequencer_csr_read -> modular_adc_0:sequencer_csr_read
	wire         mm_interconnect_0_modular_adc_0_sequencer_csr_write;        // mm_interconnect_0:modular_adc_0_sequencer_csr_write -> modular_adc_0:sequencer_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_0_sequencer_csr_writedata;    // mm_interconnect_0:modular_adc_0_sequencer_csr_writedata -> modular_adc_0:sequencer_csr_writedata
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:modular_adc_0_reset_sink_reset_bridge_in_reset_reset, modular_adc_0:reset_sink_reset_n]

	ADCTestADC_altpll_0 altpll_0 (
		.clk       (clk_clk),                        //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                               //             pll_slave.read
		.write     (),                               //                      .write
		.address   (),                               //                      .address
		.readdata  (),                               //                      .readdata
		.writedata (),                               //                      .writedata
		.c0        (altpll_0_c0_clk),                //                    c0.clk
		.locked    (altpll_0_locked_conduit_export)  //        locked_conduit.export
	);

	ADCTestADC_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	ADCTestADC_modular_adc_0 modular_adc_0 (
		.clock_clk                  (clk_clk),                                                    //            clock.clk
		.reset_sink_reset_n         (~rst_controller_reset_out_reset),                            //       reset_sink.reset_n
		.adc_pll_clock_clk          (altpll_0_c0_clk),                                            //    adc_pll_clock.clk
		.adc_pll_locked_export      (altpll_0_locked_conduit_export),                             //   adc_pll_locked.export
		.sequencer_csr_address      (mm_interconnect_0_modular_adc_0_sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (mm_interconnect_0_modular_adc_0_sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (mm_interconnect_0_modular_adc_0_sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (mm_interconnect_0_modular_adc_0_sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (mm_interconnect_0_modular_adc_0_sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (mm_interconnect_0_modular_adc_0_sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (mm_interconnect_0_modular_adc_0_sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (mm_interconnect_0_modular_adc_0_sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (mm_interconnect_0_modular_adc_0_sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (mm_interconnect_0_modular_adc_0_sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       ()                                                            // sample_store_irq.irq
	);

	ADCTestADC_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                        (clk_clk),                                                    //                                      clk_0_clk.clk
		.master_0_clk_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                             //       master_0_clk_reset_reset_bridge_in_reset.reset
		.modular_adc_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // modular_adc_0_reset_sink_reset_bridge_in_reset.reset
		.master_0_master_address                              (master_0_master_address),                                    //                                master_0_master.address
		.master_0_master_waitrequest                          (master_0_master_waitrequest),                                //                                               .waitrequest
		.master_0_master_byteenable                           (master_0_master_byteenable),                                 //                                               .byteenable
		.master_0_master_read                                 (master_0_master_read),                                       //                                               .read
		.master_0_master_readdata                             (master_0_master_readdata),                                   //                                               .readdata
		.master_0_master_readdatavalid                        (master_0_master_readdatavalid),                              //                                               .readdatavalid
		.master_0_master_write                                (master_0_master_write),                                      //                                               .write
		.master_0_master_writedata                            (master_0_master_writedata),                                  //                                               .writedata
		.modular_adc_0_sample_store_csr_address               (mm_interconnect_0_modular_adc_0_sample_store_csr_address),   //                 modular_adc_0_sample_store_csr.address
		.modular_adc_0_sample_store_csr_write                 (mm_interconnect_0_modular_adc_0_sample_store_csr_write),     //                                               .write
		.modular_adc_0_sample_store_csr_read                  (mm_interconnect_0_modular_adc_0_sample_store_csr_read),      //                                               .read
		.modular_adc_0_sample_store_csr_readdata              (mm_interconnect_0_modular_adc_0_sample_store_csr_readdata),  //                                               .readdata
		.modular_adc_0_sample_store_csr_writedata             (mm_interconnect_0_modular_adc_0_sample_store_csr_writedata), //                                               .writedata
		.modular_adc_0_sequencer_csr_address                  (mm_interconnect_0_modular_adc_0_sequencer_csr_address),      //                    modular_adc_0_sequencer_csr.address
		.modular_adc_0_sequencer_csr_write                    (mm_interconnect_0_modular_adc_0_sequencer_csr_write),        //                                               .write
		.modular_adc_0_sequencer_csr_read                     (mm_interconnect_0_modular_adc_0_sequencer_csr_read),         //                                               .read
		.modular_adc_0_sequencer_csr_readdata                 (mm_interconnect_0_modular_adc_0_sequencer_csr_readdata),     //                                               .readdata
		.modular_adc_0_sequencer_csr_writedata                (mm_interconnect_0_modular_adc_0_sequencer_csr_writedata)     //                                               .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
