//          (C) COPYRIGHT 2017 HWRACING FORMULA STUDENT TEAM
//              ALL RIGHTS RESERVED


`include "dut_if.sv"
`include "dut_wrapper.sv"
