//          (C) COPYRIGHT 2017 HWRACING FORMULA STUDENT TEAM
//              ALL RIGHTS RESERVED
// Interface for connecting the item to the DUT

interface dut_if (input clk);
  logic upBut;
  logic downBut;
  logic neturalBut;
  logic upOut;
  logic downOut;
endinterface